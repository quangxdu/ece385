library verilog;
use verilog.vl_types.all;
entity Mapper is
    port(
        DrawX           : in     vl_logic_vector(9 downto 0);
        DrawY           : in     vl_logic_vector(9 downto 0);
        PosX1           : in     vl_logic_vector(9 downto 0);
        PosY1           : in     vl_logic_vector(9 downto 0);
        PosX2           : in     vl_logic_vector(9 downto 0);
        PosY2           : in     vl_logic_vector(9 downto 0);
        PosX3           : in     vl_logic_vector(9 downto 0);
        PosY3           : in     vl_logic_vector(9 downto 0);
        PosX4           : in     vl_logic_vector(9 downto 0);
        PosY4           : in     vl_logic_vector(9 downto 0);
        PosX5           : in     vl_logic_vector(9 downto 0);
        PosY5           : in     vl_logic_vector(9 downto 0);
        PosX6           : in     vl_logic_vector(9 downto 0);
        PosY6           : in     vl_logic_vector(9 downto 0);
        PosX7           : in     vl_logic_vector(9 downto 0);
        PosY7           : in     vl_logic_vector(9 downto 0);
        PosX8           : in     vl_logic_vector(9 downto 0);
        PosY8           : in     vl_logic_vector(9 downto 0);
        PosX9           : in     vl_logic_vector(9 downto 0);
        PosY9           : in     vl_logic_vector(9 downto 0);
        PosX10          : in     vl_logic_vector(9 downto 0);
        PosY10          : in     vl_logic_vector(9 downto 0);
        PosX11          : in     vl_logic_vector(9 downto 0);
        PosY11          : in     vl_logic_vector(9 downto 0);
        PosX12          : in     vl_logic_vector(9 downto 0);
        PosY12          : in     vl_logic_vector(9 downto 0);
        PosX13          : in     vl_logic_vector(9 downto 0);
        PosY13          : in     vl_logic_vector(9 downto 0);
        PosX14          : in     vl_logic_vector(9 downto 0);
        PosY14          : in     vl_logic_vector(9 downto 0);
        PosX15          : in     vl_logic_vector(9 downto 0);
        PosY15          : in     vl_logic_vector(9 downto 0);
        PosX16          : in     vl_logic_vector(9 downto 0);
        PosY16          : in     vl_logic_vector(9 downto 0);
        SpriteID1       : in     vl_logic_vector(3 downto 0);
        SpriteID2       : in     vl_logic_vector(3 downto 0);
        SpriteID3       : in     vl_logic_vector(3 downto 0);
        SpriteID4       : in     vl_logic_vector(3 downto 0);
        SpriteID5       : in     vl_logic_vector(3 downto 0);
        SpriteID6       : in     vl_logic_vector(3 downto 0);
        SpriteID7       : in     vl_logic_vector(3 downto 0);
        SpriteID8       : in     vl_logic_vector(3 downto 0);
        SpriteID9       : in     vl_logic_vector(3 downto 0);
        SpriteID10      : in     vl_logic_vector(3 downto 0);
        SpriteID11      : in     vl_logic_vector(3 downto 0);
        SpriteID12      : in     vl_logic_vector(3 downto 0);
        SpriteID13      : in     vl_logic_vector(3 downto 0);
        SpriteID14      : in     vl_logic_vector(3 downto 0);
        SpriteID15      : in     vl_logic_vector(3 downto 0);
        SpriteID16      : in     vl_logic_vector(3 downto 0);
        spriteIDOut     : out    vl_logic_vector(3 downto 0);
        sPosXOut        : out    vl_logic_vector(4 downto 0);
        sPosYOut        : out    vl_logic_vector(4 downto 0)
    );
end Mapper;
