module GameControl
(
);

endmodule