module sprite_table(input [3:0] spriteID, input [4:0]posX, input [4:0] posY,output [7:0] color);

parameter ADDR_WIDTH = 10;
parameter DATA_WIDTH = 8;
logic [9:0] addr_reg;
parameter[0:2**10-1][7:0] Sprite0 = {
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 
8'b00000000, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000000, 
8'b00000000, 8'b00000010, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000100, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000000, 
8'b00000000, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000000, 
8'b00000000, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000110, 8'b00000110, 8'b00000100, 8'b00000000, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000100, 8'b00000000, 
8'b00000000, 8'b00000001, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000110, 8'b00000011, 8'b00000110, 8'b00000101, 8'b00000011, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000100, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000100, 8'b00000010, 8'b00001000, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00001000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00001000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000111, 8'b00000111, 8'b00000011, 8'b00001000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

	
parameter[0:2**10-1][7:0] Sprite1 = {
 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 
8'b00000000, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000000, 
8'b00000000, 8'b00000010, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000100, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000000, 
8'b00000000, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000000, 
8'b00000000, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000110, 8'b00000110, 8'b00000100, 8'b00000000, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000100, 8'b00000000, 
8'b00000000, 8'b00000001, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000110, 8'b00000011, 8'b00000110, 8'b00000101, 8'b00000011, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000100, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000100, 8'b00000010, 8'b00001000, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00001000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00001000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000111, 8'b00000111, 8'b00000011, 8'b00001000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};


parameter[0:2**10-1][7:0] Sprite2= {
 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001000, 8'b00000011, 8'b00000111, 8'b00000111, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001000, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001000, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00001000, 8'b00000010, 8'b00000100, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000100, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000011, 8'b00000101, 8'b00000110, 8'b00000011, 8'b00000110, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000001, 8'b00000000, 
8'b00000000, 8'b00000100, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000000, 8'b00000100, 8'b00000110, 8'b00000110, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000000, 
8'b00000000, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000000, 
8'b00000000, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000100, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000010, 8'b00000000, 
8'b00000000, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000000, 
8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

parameter[0:2**10-1][7:0] Sprite3= {
 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000100, 8'b00000100, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00001000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00001000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000111, 8'b00000011, 8'b00001000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00001000, 8'b00000001, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000100, 8'b00000110, 8'b00000110, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 
8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000100, 8'b00000000, 
8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000100, 8'b00000000, 
8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000110, 8'b00000100, 8'b00000111, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000111, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00000100, 8'b00000100, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

parameter[0:2**10-1][7:0] Sprite4= {
 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000100, 8'b00000100, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000001, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000111, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000111, 8'b00000100, 8'b00000110, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 
8'b00000000, 8'b00000100, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 
8'b00000000, 8'b00000100, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000000, 
8'b00000000, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000110, 8'b00000110, 8'b00000100, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000001, 8'b00001000, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001000, 8'b00000011, 8'b00000111, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001000, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001000, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00000100, 8'b00000100, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

parameter[0:2**10-1][7:0] Sprite5= {
 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000110, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00000110, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00001011, 8'b00001100, 8'b00001100, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00000010, 8'b00000010, 8'b00001100, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000110, 8'b00000110, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000001, 8'b00001100, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00000010, 8'b00000010, 8'b00001100, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00001110, 8'b00000111, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000001, 8'b00000001, 8'b00001100, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000110, 8'b00000110, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000010, 8'b00001100, 8'b00001111, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001111, 8'b00001100, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00000001, 8'b00000010, 8'b00001100, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001101, 8'b00010000, 8'b00010000, 8'b00001101, 8'b00001101, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001100, 8'b00001110, 8'b00000110, 8'b00001001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000001, 8'b00001100, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010000, 8'b00000110, 8'b00001110, 8'b00010000, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010001, 8'b00010010, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00000010, 8'b00000010, 8'b00001100, 8'b00010001, 8'b00010001, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001100, 8'b00000110, 8'b00000100, 8'b00000110, 8'b00000111, 8'b00010000, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010001, 8'b00010010, 8'b00001110, 8'b00000111, 8'b00001001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000001, 8'b00000001, 8'b00010010, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00001111, 8'b00001000, 8'b00000010, 8'b00000100, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00010000, 8'b00001111, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010010, 8'b00000110, 8'b00000110, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000010, 8'b00010011, 8'b00010100, 8'b00010100, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010101, 8'b00000001, 8'b00000001, 8'b00000111, 8'b00010010, 8'b00010010, 8'b00001010, 8'b00000110, 8'b00000111, 8'b00010000, 8'b00010100, 8'b00010100, 8'b00010001, 8'b00010001, 8'b00010100, 8'b00010010, 8'b00001110, 8'b00000111, 8'b00000111, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000111, 8'b00000001, 8'b00001011, 8'b00010010, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010001, 8'b00010110, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00010111, 8'b00001111, 8'b00001111, 8'b00010111, 8'b00001001, 8'b00000110, 8'b00000111, 8'b00001000, 8'b00010001, 8'b00010001, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010010, 8'b00000110, 8'b00000110, 8'b00001010, 8'b00000000, 
8'b00000110, 8'b00000010, 8'b00000001, 8'b00010010, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00011000, 8'b00000100, 8'b00000000, 8'b00000001, 8'b00001100, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010001, 8'b00010010, 8'b00000111, 8'b00000110, 8'b00000100, 8'b00010000, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00011001, 8'b00000110, 8'b00000111, 8'b00000110, 
8'b00000110, 8'b00000010, 8'b00000001, 8'b00010010, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010000, 8'b00001010, 8'b00000010, 8'b00000000, 8'b00000001, 8'b00010111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010001, 8'b00011010, 8'b00000111, 8'b00000110, 8'b00000010, 8'b00000010, 8'b00010101, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00011001, 8'b00001010, 8'b00001001, 8'b00000111, 
8'b00000000, 8'b00001010, 8'b00000001, 8'b00000010, 8'b00010010, 8'b00010100, 8'b00010100, 8'b00011000, 8'b00001001, 8'b00001010, 8'b00000110, 8'b00000100, 8'b00000001, 8'b00010111, 8'b00010001, 8'b00001111, 8'b00010001, 8'b00010001, 8'b00010111, 8'b00000111, 8'b00000111, 8'b00000110, 8'b00000001, 8'b00000010, 8'b00001000, 8'b00010100, 8'b00010100, 8'b00011001, 8'b00001001, 8'b00001001, 8'b00001010, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000010, 8'b00010010, 8'b00010000, 8'b00001001, 8'b00001001, 8'b00001000, 8'b00001010, 8'b00000100, 8'b00000001, 8'b00010010, 8'b00010111, 8'b00010111, 8'b00010111, 8'b00010111, 8'b00010000, 8'b00000111, 8'b00000111, 8'b00001010, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00010010, 8'b00010000, 8'b00001001, 8'b00001001, 8'b00000111, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000001, 8'b00000111, 8'b00001001, 8'b00001000, 8'b00000110, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000010, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000010, 8'b00000110, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00001010, 8'b00001001, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00000010, 8'b00000110, 8'b00001001, 8'b00000111, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00000111, 8'b00001010, 8'b00001010, 8'b00001010, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000010, 8'b00000000, 8'b00000111, 8'b00000100, 8'b00000100, 8'b00001001, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00001000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00010010, 8'b00011011, 8'b00011011, 8'b00011011, 8'b00011011, 8'b00010010, 8'b00000111, 8'b00000111, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00001000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00011010, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00011010, 8'b00001010, 8'b00001001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000100, 8'b00000001, 8'b00011100, 8'b00011101, 8'b00011101, 8'b00011101, 8'b00011101, 8'b00011100, 8'b00001001, 8'b00001001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000010, 8'b00001010, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000100, 8'b00000000, 8'b00000110, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00011110, 8'b00011111, 8'b00011011, 8'b00011011, 8'b00011111, 8'b00011001, 8'b00001001, 8'b00001001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00011110, 8'b00100000, 8'b00010100, 8'b00010100, 8'b00100000, 8'b00011110, 8'b00001001, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00011110, 8'b00011111, 8'b00011111, 8'b00011111, 8'b00011111, 8'b00100001, 8'b00001001, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000100, 8'b00000000, 8'b00000111, 8'b00001010, 8'b00001010, 8'b00001010, 8'b00001010, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00000010, 8'b00000110, 8'b00001001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

parameter[0:2**10-1][7:0] Sprite6= {
 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001000, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00000110, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001010, 8'b00001010, 8'b00001010, 8'b00001010, 8'b00000111, 8'b00000000, 8'b00000100, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00001001, 8'b00100001, 8'b00011111, 8'b00011111, 8'b00011111, 8'b00011111, 8'b00011110, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00001001, 8'b00001001, 8'b00011110, 8'b00100000, 8'b00010100, 8'b00010100, 8'b00100000, 8'b00011110, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001001, 8'b00001001, 8'b00011001, 8'b00011111, 8'b00011011, 8'b00011011, 8'b00011111, 8'b00011110, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00000110, 8'b00000000, 8'b00000100, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001010, 8'b00000010, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001001, 8'b00001001, 8'b00011100, 8'b00011101, 8'b00011101, 8'b00011101, 8'b00011101, 8'b00011100, 8'b00000001, 8'b00000100, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001001, 8'b00001010, 8'b00011010, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00011010, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00001000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000111, 8'b00000111, 8'b00010010, 8'b00011011, 8'b00011011, 8'b00011011, 8'b00011011, 8'b00010010, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00001000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00001001, 8'b00000100, 8'b00000100, 8'b00000111, 8'b00000000, 8'b00000010, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00001010, 8'b00001010, 8'b00001010, 8'b00000111, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000111, 8'b00001001, 8'b00000110, 8'b00000010, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00001001, 8'b00001010, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00000110, 8'b00000010, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000110, 8'b00000010, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000110, 8'b00001000, 8'b00001001, 8'b00000111, 8'b00000001, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000111, 8'b00001001, 8'b00001001, 8'b00010000, 8'b00010010, 8'b00000010, 8'b00000000, 8'b00000110, 8'b00001010, 8'b00000111, 8'b00000111, 8'b00010000, 8'b00010111, 8'b00010111, 8'b00010111, 8'b00010111, 8'b00010010, 8'b00000001, 8'b00000100, 8'b00001010, 8'b00001000, 8'b00001001, 8'b00001001, 8'b00010000, 8'b00010010, 8'b00000010, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00001010, 8'b00001001, 8'b00001001, 8'b00011001, 8'b00010100, 8'b00010100, 8'b00001000, 8'b00000010, 8'b00000001, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00010111, 8'b00010001, 8'b00010001, 8'b00001111, 8'b00010001, 8'b00010111, 8'b00000001, 8'b00000100, 8'b00000110, 8'b00001010, 8'b00001001, 8'b00011000, 8'b00010100, 8'b00010100, 8'b00010010, 8'b00000010, 8'b00000001, 8'b00001010, 8'b00000000, 
8'b00000111, 8'b00001001, 8'b00001010, 8'b00011001, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010101, 8'b00000010, 8'b00000010, 8'b00000110, 8'b00000111, 8'b00011010, 8'b00010001, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010111, 8'b00000001, 8'b00000000, 8'b00000010, 8'b00001010, 8'b00010000, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010010, 8'b00000001, 8'b00000010, 8'b00000110, 
8'b00000110, 8'b00000111, 8'b00000110, 8'b00011001, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010000, 8'b00000100, 8'b00000110, 8'b00000111, 8'b00010010, 8'b00010001, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001100, 8'b00000001, 8'b00000000, 8'b00000100, 8'b00011000, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010010, 8'b00000001, 8'b00000010, 8'b00000110, 
8'b00000000, 8'b00001010, 8'b00000110, 8'b00000110, 8'b00010010, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010001, 8'b00010001, 8'b00001000, 8'b00000111, 8'b00000110, 8'b00001001, 8'b00010111, 8'b00001111, 8'b00001111, 8'b00010111, 8'b00000110, 8'b00000000, 8'b00000001, 8'b00010110, 8'b00010001, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010010, 8'b00001011, 8'b00000001, 8'b00000111, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000111, 8'b00000111, 8'b00001110, 8'b00010010, 8'b00010100, 8'b00010001, 8'b00010001, 8'b00010100, 8'b00010100, 8'b00010000, 8'b00000111, 8'b00000110, 8'b00001010, 8'b00010010, 8'b00010010, 8'b00000111, 8'b00000001, 8'b00000001, 8'b00010101, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010100, 8'b00010100, 8'b00010011, 8'b00000010, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000110, 8'b00000110, 8'b00010010, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00001111, 8'b00010000, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000110, 8'b00000100, 8'b00000010, 8'b00001000, 8'b00001111, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010010, 8'b00000001, 8'b00000001, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001001, 8'b00000111, 8'b00001110, 8'b00010010, 8'b00010001, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010000, 8'b00000111, 8'b00000110, 8'b00000100, 8'b00000110, 8'b00001100, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010001, 8'b00010001, 8'b00001100, 8'b00000010, 8'b00000010, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000111, 8'b00000110, 8'b00010010, 8'b00010001, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010000, 8'b00001110, 8'b00000110, 8'b00010000, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001100, 8'b00000001, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001001, 8'b00000110, 8'b00001110, 8'b00001100, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001101, 8'b00001101, 8'b00010000, 8'b00010000, 8'b00001101, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001100, 8'b00000010, 8'b00000001, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000111, 8'b00000110, 8'b00001100, 8'b00001111, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001111, 8'b00001100, 8'b00000010, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000110, 8'b00000110, 8'b00001100, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000001, 8'b00000001, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00000111, 8'b00001110, 8'b00001100, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000010, 8'b00000010, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000111, 8'b00000110, 8'b00001100, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000001, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00000110, 8'b00000110, 8'b00001100, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000010, 8'b00000010, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00001100, 8'b00001100, 8'b00001011, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000110, 8'b00000110, 8'b00000001, 8'b00000001, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00000110, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

parameter[0:2**10-1][7:0] Sprite7= {
 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00000010, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000010, 8'b00010010, 8'b00010010, 8'b00001011, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00000010, 8'b00000010, 8'b00010010, 8'b00010100, 8'b00010100, 8'b00010010, 8'b00000010, 8'b00000001, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000001, 8'b00010010, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010011, 8'b00000001, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001000, 8'b00000110, 8'b00000111, 8'b00010000, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010010, 8'b00000010, 8'b00000010, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00011000, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010001, 8'b00001100, 8'b00000001, 8'b00000001, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00001000, 8'b00001001, 8'b00001001, 8'b00010000, 8'b00010100, 8'b00010100, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00001100, 8'b00000010, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00001000, 8'b00001010, 8'b00001010, 8'b00011000, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00001111, 8'b00001100, 8'b00000010, 8'b00000001, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00001010, 8'b00000110, 8'b00000010, 8'b00000100, 8'b00010110, 8'b00010001, 8'b00010001, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001100, 8'b00000001, 8'b00000010, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00001001, 8'b00000010, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000010, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00010101, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001100, 8'b00000010, 8'b00000010, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00001001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00001000, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000001, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00001001, 8'b00000100, 8'b00000111, 8'b00100001, 8'b00011110, 8'b00011110, 8'b00000110, 8'b00000010, 8'b00011100, 8'b00011010, 8'b00010010, 8'b00000110, 8'b00000010, 8'b00010010, 8'b00010111, 8'b00010111, 8'b00001100, 8'b00000110, 8'b00000001, 8'b00000010, 8'b00001100, 8'b00001111, 8'b00001111, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000010, 8'b00000010, 8'b00000111, 8'b00000000, 8'b00000000, 
8'b00001001, 8'b00000100, 8'b00001010, 8'b00011111, 8'b00100000, 8'b00011111, 8'b00001001, 8'b00001010, 8'b00011101, 8'b00010100, 8'b00011011, 8'b00000111, 8'b00000110, 8'b00010111, 8'b00010001, 8'b00001111, 8'b00001111, 8'b00010111, 8'b00000111, 8'b00000100, 8'b00000100, 8'b00010000, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00001011, 8'b00000001, 8'b00000111, 8'b00000000, 
8'b00001001, 8'b00000100, 8'b00001010, 8'b00011111, 8'b00010100, 8'b00011011, 8'b00001001, 8'b00001001, 8'b00011101, 8'b00010100, 8'b00011011, 8'b00001010, 8'b00000111, 8'b00010111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010010, 8'b00000110, 8'b00000100, 8'b00000110, 8'b00010000, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000001, 8'b00000010, 8'b00000110, 
8'b00001001, 8'b00000100, 8'b00001010, 8'b00011111, 8'b00010100, 8'b00011011, 8'b00001001, 8'b00001001, 8'b00011101, 8'b00010100, 8'b00011011, 8'b00001010, 8'b00000111, 8'b00010111, 8'b00010001, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00010010, 8'b00000111, 8'b00000110, 8'b00001110, 8'b00010000, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000110, 8'b00000110, 8'b00000110, 
8'b00001001, 8'b00000100, 8'b00001010, 8'b00011111, 8'b00100000, 8'b00011111, 8'b00001001, 8'b00001001, 8'b00011101, 8'b00010100, 8'b00011011, 8'b00001010, 8'b00000111, 8'b00010111, 8'b00010001, 8'b00010001, 8'b00001111, 8'b00010111, 8'b00001010, 8'b00001110, 8'b00000111, 8'b00010000, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000111, 8'b00000110, 8'b00001010, 8'b00000000, 
8'b00001001, 8'b00000010, 8'b00001001, 8'b00100001, 8'b00011110, 8'b00011001, 8'b00001001, 8'b00001001, 8'b00011100, 8'b00011010, 8'b00010010, 8'b00000111, 8'b00000111, 8'b00010000, 8'b00010111, 8'b00011010, 8'b00010010, 8'b00001001, 8'b00000110, 8'b00000111, 8'b00010000, 8'b00001111, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00000000, 8'b00000000, 
8'b00001001, 8'b00000110, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001010, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000110, 8'b00000111, 8'b00010000, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001101, 8'b00001101, 8'b00001100, 8'b00000110, 8'b00000110, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00001000, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00001001, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000111, 8'b00000110, 8'b00000110, 8'b00000111, 8'b00010000, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001100, 8'b00001110, 8'b00000111, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000010, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00001010, 8'b00000110, 8'b00000010, 8'b00000100, 8'b00001000, 8'b00010100, 8'b00010001, 8'b00001111, 8'b00001111, 8'b00001111, 8'b00001100, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000110, 8'b00000001, 8'b00000010, 8'b00010000, 8'b00010001, 8'b00010100, 8'b00010001, 8'b00001111, 8'b00010001, 8'b00001100, 8'b00000110, 8'b00000110, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000110, 8'b00000000, 8'b00000010, 8'b00010101, 8'b00010100, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010001, 8'b00010010, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000110, 8'b00000100, 8'b00000001, 8'b00000010, 8'b00001000, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010001, 8'b00010010, 8'b00000110, 8'b00000110, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00001000, 8'b00000100, 8'b00000110, 8'b00010010, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010010, 8'b00001110, 8'b00000111, 8'b00001001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00001001, 8'b00001010, 8'b00010000, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010100, 8'b00010010, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00001001, 8'b00001001, 8'b00011001, 8'b00010100, 8'b00010100, 8'b00010010, 8'b00001110, 8'b00000110, 8'b00001001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00001001, 8'b00001001, 8'b00011001, 8'b00011001, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00001001, 8'b00001010, 8'b00000110, 8'b00000110, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001010, 8'b00001001, 8'b00000111, 8'b00001010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

parameter[0:2**10-1][7:0] Sprite15= {
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

parameter[0:2**10-1][7:0] Sprite8= {
 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001011, 8'b00100010, 8'b00100010, 8'b00100011, 8'b00100010, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00100010, 8'b00100010, 8'b00100010, 8'b00100100, 8'b00100010, 8'b00100010, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100100, 8'b00100010, 8'b00100100, 8'b00100100, 8'b00100100, 8'b00100010, 8'b00100010, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100010, 8'b00100010, 8'b00100101, 8'b00100100, 8'b00100100, 8'b00100010, 8'b00100011, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100010, 8'b00100010, 8'b00100101, 8'b00100100, 8'b00100100, 8'b00100010, 8'b00100011, 8'b00100101, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100010, 8'b00100010, 8'b00001011, 8'b00100100, 8'b00100100, 8'b00100100, 8'b00100011, 8'b00001011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100100, 8'b00100010, 8'b00001011, 8'b00100100, 8'b00100100, 8'b00100100, 8'b00100010, 8'b00100100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100100, 8'b00100011, 8'b00100100, 8'b00100100, 8'b00100010, 8'b00100100, 8'b00100010, 8'b00100010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001011, 8'b00100011, 8'b00100100, 8'b00100100, 8'b00100010, 8'b00100100, 8'b00100010, 8'b00100011, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100011, 8'b00100100, 8'b00100100, 8'b00100010, 8'b00100010, 8'b00100010, 8'b00100011, 8'b00100010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100010, 8'b00100010, 8'b00100100, 8'b00100010, 8'b00100010, 8'b00100010, 8'b00100010, 8'b00100011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001011, 8'b00100011, 8'b00100100, 8'b00100010, 8'b00100010, 8'b00100010, 8'b00100010, 8'b00100011, 8'b00001011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100011, 8'b00100100, 8'b00100010, 8'b00100110, 8'b00100110, 8'b00100010, 8'b00100010, 8'b00100011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100101, 8'b00100011, 8'b00100011, 8'b00100101, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100010, 8'b00100010, 8'b00100010, 8'b00100110, 8'b00100110, 8'b00100110, 8'b00100010, 8'b00100011, 8'b00001011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100011, 8'b00100010, 8'b00100010, 8'b00100011, 8'b00100100, 8'b00000000, 8'b00000000, 8'b00001011, 8'b00100011, 8'b00100100, 8'b00100110, 8'b00100110, 8'b00100110, 8'b00100010, 8'b00100010, 8'b00100011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100011, 8'b00100010, 8'b00100010, 8'b00100010, 8'b00100100, 8'b00100011, 8'b00100010, 8'b00000000, 8'b00100011, 8'b00100010, 8'b00100010, 8'b00100111, 8'b00100111, 8'b00100011, 8'b00100010, 8'b00100011, 8'b00100100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100011, 8'b00100010, 8'b00100010, 8'b00100111, 8'b00100111, 8'b00100010, 8'b00100100, 8'b00100011, 8'b00101000, 8'b00100011, 8'b00100010, 8'b00100111, 8'b00100111, 8'b00100111, 8'b00100011, 8'b00100010, 8'b00100011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00100011, 8'b00100010, 8'b00100010, 8'b00100111, 8'b00100111, 8'b00100111, 8'b00100111, 8'b00100011, 8'b00100010, 8'b00100010, 8'b00100010, 8'b00100011, 8'b00100111, 8'b00100111, 8'b00100111, 8'b00100011, 8'b00100011, 8'b00100010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00101000, 8'b00100011, 8'b00100011, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00100010, 8'b00100011, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00100011, 8'b00101000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00001011, 8'b00101000, 8'b00100011, 8'b00100111, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101001, 8'b00101000, 8'b00100011, 8'b00100011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001011, 8'b00101000, 8'b00101000, 8'b00101000, 8'b00101001, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101000, 8'b00101000, 8'b00100100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001011, 8'b00101011, 8'b00101000, 8'b00101001, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101000, 8'b00101011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001011, 8'b00101011, 8'b00101000, 8'b00101000, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101010, 8'b00101000, 8'b00101000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001011, 8'b00101011, 8'b00101000, 8'b00101001, 8'b00101010, 8'b00101100, 8'b00101100, 8'b00101100, 8'b00101100, 8'b00101011, 8'b00101011, 8'b00100010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001011, 8'b00101011, 8'b00000110, 8'b00101011, 8'b00101011, 8'b00101011, 8'b00101011, 8'b00101011, 8'b00101011, 8'b00101101, 8'b00100100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000011, 8'b00011010, 8'b00011010, 8'b00011010, 8'b00011010, 8'b00011010, 8'b00011010, 8'b00011010, 8'b00101101, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
};
parameter[0:2**10-1][7:0] Sprite9= {
 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101110, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00101110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00110000, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00110000, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00110000, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00110000, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110000, 8'b00000000, 
8'b00101110, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00101110, 
8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00001011, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 
8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00001011, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 8'b00000000, 
8'b00101111, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00101111, 
8'b00101110, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00101110, 
8'b00000000, 8'b00110000, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00110000, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00110000, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110001, 8'b00110001, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00110000, 8'b00110001, 8'b00110010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00110010, 8'b00110001, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101110, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00101110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
};


logic [7:0]sprite0color;
logic [7:0]sprite1color;
logic [7:0]sprite2color;
logic [7:0]sprite3color;
logic [7:0]sprite4color;
logic [7:0]sprite5color;
logic [7:0]sprite6color;
logic [7:0]sprite7color;
logic [7:0]sprite8color;
logic [7:0]sprite9color;
logic [7:0]sprite15color;
assign sprite15color=Sprite15[(32*int'(posY)+int'(posX))];
assign sprite0color=Sprite0[(32*int'(posY)+int'(posX))];
assign sprite1color=Sprite1[(32*int'(posY)+int'(posX))];
assign sprite2color=Sprite2[(32*int'(posY)+int'(posX))];
assign sprite3color=Sprite3[(32*int'(posY)+int'(posX))];
assign sprite4color=Sprite4[(32*int'(posY)+int'(posX))];
assign sprite5color=Sprite5[(32*int'(posY)+int'(posX))];
assign sprite6color=Sprite6[(32*int'(posY)+int'(posX))];
assign sprite7color=Sprite7[(32*int'(posY)+int'(posX))];
assign sprite8color=Sprite8[(32*int'(posY)+int'(posX))];
assign sprite9color=Sprite9[(32*int'(posY)+int'(posX))];

mux16 mux16
(
	.sel(spriteID),
	.i1(sprite0color),
	.i2(sprite1color),
	.i3(sprite2color),
	.i4(sprite3color),
	.i5(sprite4color),
	.i6(sprite5color),
	.i7(sprite6color),
	.i8(sprite7color),
	.i9(sprite8color),
	.i10(sprite9color),
	.i11(sprite15color),
	.i12(sprite15color),
	.i13(sprite15color),
	.i14(sprite15color),
	.i15(sprite15color),
	.i16(sprite15color),
	.f(color)
);

endmodule
